//***************************************************************************//
//***************************************************************************//
//***************************************************************************//
//**************                                          *******************//
//**************                                          *******************//
//**************      (c) SASIC Technologies Pvt Ltd      *******************//
//**************          (c) Verilogic Solutions         *******************//
//**************                                          *******************//
//**************                                          *******************//
//**************                                          *******************//
//**************           www.sasictek.com               *******************//
//**************          www.verilog-ic.com              *******************//
//**************                                          *******************//
//**************           Twitter:@sasictek              *******************//
//**************                                          *******************//
//**************                                          *******************//
//**************                                          *******************//
//***************************************************************************//
//***************************************************************************//


//              File Name : apb.interface.sv
//              File Type: System Verilog                                 
//              Creation Date : 22-02-2017
//              Last Modified : Tue 28 Feb 2017 02:42:39 PM IST

                             
//***************************************************************************//
//***************************************************************************//
                             

//              Author:
//              Reviewer:
//              Manager:
                             

//***************************************************************************//
//***************************************************************************//

//import apb_package::*;

interface apb_interface(input logic top_clk);

logic prst;
logic psel;
logic penable;
logic pwr;
logic [ADD_WIDTH-1:0]padd;
logic [DATA_WIDTH-1:0]pwdata;
logic [DATA_WIDTH-1:0]prdata;
logic pslverr;
logic pready;

clocking drv_cb@(negedge top_clk);

	output prst;
	output psel;
	output penable;
	output pwr;
	output padd;
	output pwdata;
	input prdata;
	input pslverr;
	input pready;
//	input top_clk;
	
	endclocking

endinterface

