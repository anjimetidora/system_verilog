//***************************************************************************//
//***************************************************************************//
//***************************************************************************//
//**************                                          *******************//
//**************                                          *******************//
//**************      (c) SASIC Technologies Pvt Ltd      *******************//
//**************          (c) Verilogic Solutions         *******************//
//**************                                          *******************//
//**************                                          *******************//
//**************                                          *******************//
//**************           www.sasictek.com               *******************//
//**************          www.verilog-ic.com              *******************//
//**************                                          *******************//
//**************           Twitter:@sasictek              *******************//
//**************                                          *******************//
//**************                                          *******************//
//**************                                          *******************//
//***************************************************************************//
//***************************************************************************//


//              File Name :                                 
//              File Type: System Verilog                                 
//              Creation Date : 20-02-2017
//              Last Modified : Fri 03 Mar 2017 11:40:37 AM IST

                             
//***************************************************************************//
//***************************************************************************//
                             

//              Author:
//              Reviewer:
//              Manager:
                             

//***************************************************************************//
//***************************************************************************//
import apb_package::*;
typedef enum bit[1:0]{READ,WRITE,RST}op;

class apb_transaction;
	logic pclk;
	logic prst;
	logic psel;
	logic penable;
	logic pwr;
	randc op kind;
	rand logic [ADD_WIDTH-1:0]padd;	//address width 4 bits
	randc logic [DATA_WIDTH-1:0]pwdata;	//data width 32 bits
	logic [DATA_WIDTH-1:0]prdata;
	logic  pslverr;
	logic  pready;

	constraint c_add{
										padd<25;
									}

	constraint c_wdata{
											pwdata>0;
											pwdata<100;}
endclass
