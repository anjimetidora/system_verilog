//***************************************************************************//
//***************************************************************************//
//***************************************************************************//
//**************                                          *******************//
//**************                                          *******************//
//**************      (c) SASIC Technologies Pvt Ltd      *******************//
//**************          (c) Verilogic Solutions         *******************//
//**************                                          *******************//
//**************                                          *******************//
//**************                                          *******************//
//**************           www.sasictek.com               *******************//
//**************          www.verilog-ic.com              *******************//
//**************                                          *******************//
//**************           Twitter:@sasictek              *******************//
//**************                                          *******************//
//**************                                          *******************//
//**************                                          *******************//
//***************************************************************************//
//***************************************************************************//


//              File Name : apb_top.sv
//              File Type: System Verilog                                 
//              Creation Date : 22-02-2017
//              Last Modified : Fri 28 Jul 2017 09:04:45 PM IST

                             
//***************************************************************************//
//***************************************************************************//
                             

//              Author:
//              Reviewer:
//              Manager:
                             

//***************************************************************************//
//***************************************************************************//

import apb_package::*;
`include"apb_environment.sv"

module apb_top;
logic top_clk;

apb_interface top_inf(.top_clk(top_clk));

apb_slave dut_insta(.*,	
							.pclk(top_clk),
              .prst(top_inf.prst),
							.psel(top_inf.psel),
							.penable(top_inf.penable),
							.pwr(top_inf.pwr),
							.padd(top_inf.padd),
							.pwdata(top_inf.pwdata),
							.prdata(top_inf.prdata),
							.pslverr(top_inf.pslverr),
							.pready(top_inf.pready)
							);

apb_environment top_env;

initial begin
top_clk='b0;
forever #5 top_clk=~top_clk;
end

initial begin
top_env=new(top_inf);
top_env.main();
#10;
$finish;
end
endmodule



